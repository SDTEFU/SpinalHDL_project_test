// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : template
// Git hash  : a62e70eb2f73b048f5ccdee8b8fff3a499db741e

`timescale 1ns/1ps

module template (
);



endmodule
