// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : template

`timescale 1ns/1ps

module template (
  input               io_inin,
  output              io_outout
);


  assign io_outout = io_inin;

endmodule
