// Generator : SpinalHDL v1.8.1    git head : 2a7592004363e5b40ec43e1f122ed8641cd8965b
// Component : template
// Git hash  : e00b864ca882cd5051405ee12ee645eec6f513e2

`timescale 1ns/1ps

module template (
);



endmodule
